`timescale 1ns / 1ps

module num_to_coins(
    input wire [8:0] number,
    output wire [13:0] value
    );

//

endmodule