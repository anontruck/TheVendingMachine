`timescale 1ns / 1ps

module num_to_7SD(
    input wire [13:0] number,
    input wire decimal,
    output wire [31:0] display
    );

//

endmodule